.SUBCKT test_passives TheBigNode

R1 TheBigNode 0
C1 TheBigNode 0
L1 TheBigNode 0

.ENDS

