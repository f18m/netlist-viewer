.SUBCKT test_passives TheBigNode

R1 TheBigNode 0 1k
C1 TheBigNode 0 1p
L1 TheBigNode 0 1u

.ENDS

